// design_under_test.sv
module design_module_name ();  // Design under test
  initial $display("Hello from design!");  // Display message
endmodule